// Creates the 64x32:1 mux.

`timescale 10ps/1ps
module big_daddy_elon_mux (
input logic [31:0][63:0] input_data,
output logic [63:0] output_data,
input logic [4:0] selects
);

	genvar i, j;
	
	logic [31:0] temp_var [63:0];
	generate
		for (i = 63; i >= 0; i--) begin: muxes
			for (j = 31; j >= 0; j--) begin: registers
				assign temp_var[i][j] = input_data[j][i];
			end
			
			mux32_1 mux_i(.out(output_data[i]), .inputs(temp_var[i]), .select(selects)); // Combines 64 32:1 muxes to create a 64x32:1 mux.
		end
	endgenerate
endmodule

module big_daddy_elon_mux_testbench();  // tests all possible select variations with an alternating input.
  logic  [31:0][63:0] input_data;
  logic  [63:0] output_data;  
  logic  [4:0] selects;      
       
  big_daddy_elon_mux dut (.input_data, .output_data, .selects);      
     
  integer i;   
  initial begin   
	 input_data[0] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[1] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[2] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[3] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[4] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[5] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[6] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[7] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[8] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[9] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[10] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[11] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[12] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[13] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[14] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[15] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[16] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[17] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[18] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[19] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[20] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[21] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[22] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[23] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[24] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[25] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[26] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[27] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[28] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[29] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	 input_data[30] = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	 input_data[31] = 64'b0000000000000000000000000000000000000000000000000000000000000000; #(960);
    
	 for(i=0; i< 32; i++) begin   
      {selects} = i; #30;    
    end   
  end   
endmodule



